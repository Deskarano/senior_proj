library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity main_tb is
--  Port ( );
end main_tb;

architecture Behavioral of main_tb is
    component main
        port( 
                clk         : in std_logic;
                int_btn     : in std_logic_vector(3 downto 0);
                leds        : out std_logic_vector(3 downto 0);
                uart_rx_pin : in std_logic;
                uart_tx_pin : out std_logic
             );
    end component;
    
    component uart_tx6
        port (
                data_in             : in std_logic_vector(7 downto 0);
                en_16_x_baud        : in std_logic;
                serial_out          : out std_logic;
                buffer_write        : in std_logic;
                buffer_data_present : out std_logic;
                buffer_half_full    : out std_logic;
                buffer_full         : out std_logic;
                buffer_reset        : in std_logic;
                clk                 : in std_logic);
    end component;
    
    component uart_rx6
        port (
                serial_in           : in std_logic;
                en_16_x_baud        : in std_logic;
                data_out            : out std_logic_vector(7 downto 0);
                buffer_read         : in std_logic;
                buffer_data_present : out std_logic;
                buffer_half_full    : out std_logic;
                buffer_full         : out std_logic;
                buffer_reset        : in std_logic;
                clk                 : in std_logic);
    end component;
    
    component sim_clk_wrapper
        port (
                sim_clk_out : out std_logic;
                sim_rst_out : out std_logic
            );
    end component;
    
    signal clk_sig : std_logic;
    signal rst_sig : std_logic;
    
    signal main_uart_rx : std_logic;
    signal main_uart_tx : std_logic;
    
    -- stuff for the UART
    signal uart_baud_count   : integer range 0 to 53        := 0;
    signal uart_baud         : std_logic                    := '0';

    signal uart_tx_buf_pres  : std_logic                    := '0';
    signal uart_tx_buf_half  : std_logic                    := '0';
    signal uart_tx_buf_full  : std_logic                    := '0';
    signal uart_rx_buf_pres  : std_logic                    := '0';
    signal uart_rx_buf_half  : std_logic                    := '0';
    signal uart_rx_buf_full  : std_logic                    := '0';
    signal uart_data_in      : std_logic_vector(7 downto 0) := (others => '0');
    signal uart_data_out     : std_logic_vector(7 downto 0) := (others => '0');
    signal uart_buffer_write : std_logic                    := '0';
    signal uart_buffer_read  : std_logic                    := '0';
    signal uart_reset        : std_logic                    := '0';
    
    -- main signals
    signal main_int_btn      : std_logic_vector(3 downto 0) := (others => '0');
    signal main_leds         : std_logic_vector(3 downto 0) := (others => '0');
begin
    sim_clk_gen : sim_clk_wrapper
        port map(
                    sim_clk_out => clk_sig,
                    sim_rst_out => rst_sig
                );
                
    sim_uart_tx : uart_tx6
        port map (
                    data_in             => uart_data_in,
                    en_16_x_baud        => uart_baud,
                    serial_out          => main_uart_rx,
                    buffer_write        => uart_buffer_write,
                    buffer_data_present => uart_tx_buf_pres,
                    buffer_half_full    => uart_tx_buf_half,
                    buffer_full         => uart_tx_buf_full,
                    buffer_reset        => uart_reset,
                    clk                 => clk_sig);
                    
    sim_uart_rx : uart_rx6
        port map ( 
                    serial_in           => main_uart_tx,
                    en_16_x_baud        => uart_baud,
                    data_out            => uart_data_out,
                    buffer_read         => uart_buffer_read,
                    buffer_data_present => uart_rx_buf_pres,
                    buffer_half_full    => uart_rx_buf_half,
                    buffer_full         => uart_rx_buf_full,
                    buffer_reset        => uart_reset,
                    clk                 => clk_sig);

    UUT : main
        port map ( 
                    clk         => clk_sig,
                    int_btn     => main_int_btn,
                    leds        => main_leds,
                    uart_rx_pin => main_uart_rx,
                    uart_tx_pin => main_uart_tx
                  );

    baud_rate: process(clk_sig)
    begin
        if rising_edge(clk_sig) then
            if uart_baud_count = 53 then
                uart_baud_count <= 0;
                uart_baud <= '1';
            else
                uart_baud_count <= uart_baud_count + 1;
                uart_baud <= '0';
            end if;
        end if;
    end process baud_rate;
    
    simulate: process
    begin
        wait for 1000us;
        wait until rising_edge(clk_sig);
        -- trigger an interrupt
        main_int_btn(0) <= '1';
        
        wait until rising_edge(clk_sig);
        wait until rising_edge(clk_sig);
        
        main_int_btn(0) <= '0';       
        uart_buffer_write <= '1';
        
        -- length
        uart_buffer_write <= '1';
        uart_data_in <= x"d4";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"07";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 0
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"10";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"11";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 2
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"12";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 3
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"13";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 4
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"14";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 5
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"15";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 6
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"16";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 7
        uart_buffer_write <= '1';
        uart_data_in <= x"01";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"80";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"02";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 8
        uart_buffer_write <= '1';
        uart_data_in <= x"04";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"d6";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"02";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 9
        uart_buffer_write <= '1';
        uart_data_in <= x"0f";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"02";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 10
        uart_buffer_write <= '1';
        uart_data_in <= x"01";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"16";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"01";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 11
        uart_buffer_write <= '1';
        uart_data_in <= x"10";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"d6";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"01";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 12
        uart_buffer_write <= '1';
        uart_data_in <= x"08";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"60";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"03";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 13
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"16";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 14
        uart_buffer_write <= '1';
        uart_data_in <= x"08";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"20";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"02";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 15
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"17";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 16
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"18";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 17
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"19";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 18
        uart_buffer_write <= '1';
        uart_data_in <= x"01";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"17";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"01";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 19
        uart_buffer_write <= '1';
        uart_data_in <= x"ff";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"d7";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"01";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 20
        uart_buffer_write <= '1';
        uart_data_in <= x"12";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"60";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"03";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 21
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"17";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 22
        uart_buffer_write <= '1';
        uart_data_in <= x"01";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"18";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"01";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 23
        uart_buffer_write <= '1';
        uart_data_in <= x"ff";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"d8";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"01";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 24
        uart_buffer_write <= '1';
        uart_data_in <= x"12";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"60";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"03";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 25
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"17";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 26
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"18";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 27
        uart_buffer_write <= '1';
        uart_data_in <= x"01";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"19";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"01";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 28
        uart_buffer_write <= '1';
        uart_data_in <= x"ff";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"d9";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"01";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 29
        uart_buffer_write <= '1';
        uart_data_in <= x"12";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"60";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"03";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 30
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"17";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 31
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"18";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 32
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"19";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 33
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"50";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"02";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 34
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 35
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 36
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 37
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 38
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 39
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 40
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 41
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 42
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 43
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 44
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 45
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 46
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 47
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 48
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 49
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 50
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 51
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 52
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 53
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 54
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 55
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 56
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 57
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 58
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 59
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 60
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 61
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 62
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 63
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 64
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 65
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 66
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 67
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 68
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 69
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 70
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 71
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 72
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 73
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 74
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 75
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 76
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 77
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 78
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 79
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 80
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 81
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 82
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 83
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 84
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 85
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 86
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 87
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 88
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 89
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 90
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 91
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 92
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 93
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 94
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 95
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 96
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 97
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 98
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 99
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 100
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 101
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 102
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 103
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 104
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 105
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 106
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 107
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 108
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 109
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 110
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 111
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 112
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 113
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 114
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 115
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 116
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 117
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 118
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 119
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 120
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 121
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 122
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 123
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 124
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 125
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 126
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 127
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 128
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 129
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 130
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 131
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 132
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 133
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 134
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 135
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 136
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 137
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 138
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 139
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 140
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 141
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 142
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 143
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 144
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 145
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 146
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 147
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 148
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 149
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 150
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 151
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 152
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 153
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 154
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 155
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 156
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 157
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 158
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 159
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 160
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 161
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 162
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 163
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 164
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 165
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 166
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 167
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 168
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 169
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 170
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 171
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 172
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 173
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 174
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 175
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 176
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 177
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 178
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 179
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 180
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 181
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 182
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 183
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 184
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 185
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 186
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 187
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 188
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 189
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 190
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 191
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 192
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 193
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 194
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 195
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 196
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 197
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 198
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 199
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 200
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 201
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 202
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 203
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 204
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 205
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 206
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 207
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 208
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 209
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 210
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 211
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 212
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 213
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 214
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 215
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 216
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 217
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 218
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 219
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 220
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 221
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 222
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 223
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 224
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 225
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 226
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 227
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 228
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 229
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 230
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 231
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 232
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 233
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 234
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 235
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 236
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 237
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 238
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 239
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 240
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 241
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 242
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 243
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 244
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 245
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 246
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 247
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 248
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 249
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 250
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 251
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 252
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 253
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 254
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 255
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 256
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 257
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 258
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 259
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 260
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 261
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 262
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 263
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 264
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 265
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 266
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 267
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 268
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 269
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 270
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 271
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 272
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 273
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 274
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 275
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 276
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 277
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 278
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 279
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 280
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 281
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 282
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 283
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 284
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 285
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 286
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 287
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 288
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 289
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 290
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 291
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 292
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 293
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 294
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 295
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 296
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 297
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 298
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 299
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 300
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 301
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 302
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 303
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 304
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 305
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 306
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 307
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 308
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 309
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 310
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 311
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 312
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 313
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 314
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 315
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 316
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 317
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 318
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 319
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 320
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 321
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 322
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 323
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 324
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 325
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 326
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 327
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 328
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 329
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 330
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 331
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 332
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 333
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 334
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 335
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 336
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 337
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 338
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 339
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 340
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 341
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 342
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 343
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 344
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 345
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 346
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 347
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 348
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 349
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 350
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 351
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 352
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 353
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 354
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 355
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 356
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 357
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 358
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 359
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 360
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 361
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 362
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 363
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 364
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 365
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 366
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 367
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 368
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 369
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 370
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 371
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 372
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 373
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 374
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 375
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 376
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 377
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 378
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 379
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 380
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 381
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 382
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 383
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 384
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 385
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 386
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 387
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 388
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 389
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 390
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 391
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 392
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 393
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 394
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 395
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 396
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 397
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 398
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 399
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 400
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 401
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 402
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 403
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 404
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 405
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 406
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 407
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 408
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 409
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 410
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 411
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 412
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 413
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 414
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 415
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 416
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 417
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 418
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 419
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 420
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 421
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 422
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 423
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 424
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 425
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 426
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 427
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 428
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 429
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 430
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 431
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 432
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 433
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 434
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 435
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 436
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 437
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 438
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 439
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 440
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 441
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 442
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 443
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 444
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 445
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 446
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 447
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 448
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 449
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 450
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 451
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 452
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 453
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 454
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 455
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 456
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 457
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 458
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 459
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 460
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 461
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 462
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 463
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 464
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 465
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 466
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 467
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 468
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 469
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 470
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 471
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 472
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 473
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 474
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 475
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 476
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 477
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 478
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 479
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 480
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 481
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 482
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 483
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 484
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 485
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 486
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 487
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 488
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 489
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 490
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 491
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 492
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 493
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 494
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 495
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 496
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 497
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 498
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 499
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 500
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 501
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 502
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 503
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 504
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 505
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 506
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 507
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 508
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 509
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 510
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 511
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 512
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 513
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 514
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 515
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 516
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 517
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 518
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 519
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 520
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 521
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 522
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 523
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 524
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 525
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 526
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 527
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 528
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 529
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 530
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 531
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 532
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 533
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 534
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 535
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 536
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 537
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 538
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 539
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 540
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 541
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 542
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 543
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 544
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 545
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 546
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 547
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 548
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 549
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 550
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 551
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 552
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 553
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 554
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 555
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 556
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 557
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 558
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 559
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 560
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 561
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 562
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 563
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 564
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 565
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 566
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 567
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 568
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 569
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 570
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 571
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 572
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 573
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 574
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 575
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 576
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 577
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 578
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 579
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 580
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 581
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 582
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 583
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 584
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 585
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 586
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 587
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 588
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 589
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 590
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 591
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 592
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 593
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 594
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 595
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 596
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 597
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 598
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 599
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 600
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 601
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 602
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 603
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 604
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 605
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 606
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 607
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 608
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 609
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 610
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 611
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 612
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 613
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 614
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 615
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 616
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 617
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 618
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 619
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 620
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 621
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 622
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 623
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 624
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 625
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 626
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 627
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 628
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 629
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 630
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 631
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 632
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 633
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 634
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 635
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 636
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 637
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 638
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 639
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 640
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 641
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 642
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 643
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 644
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 645
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 646
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 647
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 648
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 649
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 650
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 651
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 652
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 653
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 654
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 655
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 656
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 657
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 658
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 659
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 660
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 661
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 662
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 663
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 664
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 665
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 666
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 667
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 668
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 669
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 670
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 671
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 672
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 673
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 674
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 675
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 676
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 677
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 678
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 679
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 680
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 681
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 682
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 683
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 684
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 685
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 686
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 687
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 688
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 689
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 690
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 691
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 692
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 693
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 694
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 695
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 696
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 697
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 698
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 699
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 700
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 701
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 702
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 703
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 704
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 705
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 706
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 707
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 708
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 709
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 710
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 711
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 712
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 713
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 714
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 715
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 716
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 717
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 718
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 719
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 720
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 721
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 722
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 723
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 724
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 725
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 726
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 727
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 728
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 729
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 730
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 731
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 732
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 733
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 734
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 735
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 736
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 737
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 738
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 739
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 740
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 741
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 742
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 743
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 744
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 745
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 746
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 747
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 748
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 749
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 750
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 751
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 752
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 753
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 754
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 755
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 756
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 757
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 758
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 759
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 760
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 761
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 762
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 763
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 764
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 765
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 766
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 767
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 768
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 769
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 770
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 771
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 772
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 773
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 774
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 775
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 776
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 777
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 778
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 779
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 780
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 781
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 782
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 783
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 784
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 785
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 786
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 787
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 788
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 789
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 790
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 791
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 792
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 793
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 794
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 795
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 796
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 797
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 798
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 799
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 800
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 801
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 802
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 803
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 804
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 805
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 806
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 807
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 808
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 809
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 810
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 811
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 812
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 813
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 814
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 815
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 816
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 817
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 818
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 819
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 820
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 821
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 822
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 823
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 824
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 825
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 826
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 827
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 828
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 829
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 830
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 831
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 832
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 833
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 834
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 835
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 836
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 837
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 838
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 839
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 840
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 841
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 842
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 843
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 844
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 845
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 846
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 847
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 848
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 849
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 850
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 851
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 852
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 853
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 854
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 855
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 856
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 857
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 858
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 859
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 860
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 861
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 862
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 863
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 864
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 865
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 866
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 867
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 868
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 869
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 870
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 871
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 872
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 873
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 874
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 875
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 876
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 877
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 878
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 879
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 880
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 881
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 882
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 883
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 884
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 885
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 886
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 887
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 888
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 889
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 890
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 891
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 892
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 893
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 894
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 895
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 896
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 897
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 898
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 899
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 900
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 901
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 902
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 903
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 904
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 905
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 906
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 907
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 908
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 909
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 910
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 911
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 912
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 913
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 914
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 915
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 916
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 917
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 918
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 919
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 920
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 921
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 922
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 923
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 924
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 925
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 926
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 927
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 928
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 929
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 930
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 931
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 932
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 933
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 934
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 935
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 936
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 937
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 938
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 939
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 940
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 941
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 942
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 943
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 944
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 945
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 946
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 947
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 948
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 949
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 950
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 951
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 952
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 953
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 954
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 955
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 956
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 957
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 958
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 959
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 960
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 961
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 962
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 963
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 964
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 965
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 966
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 967
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 968
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 969
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 970
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 971
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 972
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 973
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 974
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 975
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 976
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 977
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 978
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 979
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 980
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 981
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 982
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 983
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 984
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 985
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 986
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 987
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 988
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 989
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 990
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 991
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 992
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 993
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 994
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 995
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 996
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 997
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 998
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 999
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1000
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1001
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1002
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1003
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1004
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1005
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1006
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1007
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1008
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1009
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1010
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1011
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1012
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1013
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1014
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1015
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1016
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1017
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1018
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1019
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1020
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1021
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1022
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1023
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1024
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1025
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1026
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1027
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1028
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1029
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1030
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1031
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1032
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1033
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1034
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1035
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1036
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1037
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1038
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1039
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1040
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1041
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1042
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1043
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1044
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1045
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1046
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1047
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1048
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1049
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1050
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1051
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1052
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1053
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1054
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1055
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1056
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1057
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1058
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1059
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1060
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1061
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1062
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1063
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1064
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1065
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1066
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1067
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1068
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1069
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1070
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1071
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1072
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1073
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1074
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1075
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1076
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1077
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1078
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1079
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1080
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1081
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1082
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1083
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1084
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1085
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1086
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1087
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1088
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1089
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1090
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1091
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1092
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1093
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1094
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1095
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1096
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1097
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1098
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1099
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1100
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1101
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1102
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1103
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1104
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1105
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1106
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1107
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1108
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1109
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1110
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1111
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1112
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1113
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1114
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1115
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1116
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1117
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1118
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1119
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1120
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1121
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1122
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1123
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1124
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1125
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1126
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1127
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1128
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1129
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1130
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1131
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1132
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1133
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1134
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1135
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1136
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1137
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1138
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1139
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1140
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1141
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1142
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1143
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1144
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1145
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1146
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1147
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1148
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1149
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1150
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1151
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1152
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1153
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1154
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1155
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1156
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1157
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1158
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1159
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1160
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1161
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1162
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1163
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1164
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1165
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1166
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1167
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1168
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1169
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1170
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1171
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1172
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1173
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1174
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1175
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1176
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1177
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1178
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1179
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1180
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1181
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1182
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1183
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1184
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1185
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1186
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1187
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1188
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1189
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1190
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1191
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1192
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1193
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1194
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1195
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1196
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1197
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1198
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1199
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1200
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1201
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1202
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1203
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1204
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1205
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1206
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1207
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1208
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1209
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1210
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1211
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1212
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1213
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1214
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1215
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1216
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1217
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1218
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1219
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1220
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1221
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1222
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1223
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1224
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1225
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1226
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1227
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1228
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1229
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1230
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1231
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1232
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1233
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1234
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1235
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1236
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1237
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1238
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1239
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1240
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1241
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1242
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1243
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1244
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1245
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1246
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1247
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1248
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1249
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1250
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1251
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1252
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1253
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1254
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1255
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1256
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1257
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1258
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1259
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1260
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1261
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1262
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1263
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1264
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1265
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1266
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1267
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1268
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1269
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1270
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1271
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1272
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1273
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1274
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1275
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1276
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1277
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1278
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1279
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1280
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1281
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1282
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1283
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1284
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1285
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1286
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1287
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1288
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1289
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1290
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1291
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1292
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1293
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1294
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1295
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1296
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1297
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1298
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1299
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1300
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1301
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1302
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1303
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1304
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1305
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1306
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1307
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1308
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1309
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1310
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1311
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1312
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1313
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1314
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1315
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1316
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1317
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1318
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1319
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1320
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1321
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1322
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1323
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1324
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1325
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1326
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1327
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1328
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1329
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1330
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1331
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1332
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1333
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1334
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1335
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1336
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1337
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1338
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1339
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1340
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1341
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1342
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1343
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1344
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1345
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1346
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1347
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1348
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1349
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1350
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1351
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1352
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1353
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1354
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1355
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1356
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1357
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1358
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1359
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1360
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1361
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1362
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1363
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1364
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1365
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1366
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1367
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1368
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1369
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1370
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1371
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1372
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1373
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1374
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1375
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1376
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1377
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1378
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1379
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1380
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1381
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1382
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1383
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1384
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1385
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1386
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1387
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1388
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1389
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1390
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1391
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1392
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1393
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1394
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1395
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1396
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1397
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1398
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1399
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1400
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1401
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1402
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1403
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1404
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1405
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1406
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1407
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1408
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1409
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1410
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1411
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1412
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1413
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1414
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1415
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1416
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1417
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1418
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1419
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1420
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1421
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1422
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1423
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1424
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1425
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1426
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1427
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1428
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1429
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1430
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1431
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1432
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1433
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1434
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1435
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1436
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1437
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1438
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1439
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1440
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1441
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1442
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1443
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1444
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1445
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1446
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1447
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1448
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1449
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1450
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1451
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1452
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1453
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1454
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1455
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1456
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1457
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1458
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1459
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1460
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1461
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1462
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1463
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1464
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1465
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1466
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1467
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1468
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1469
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1470
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1471
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1472
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1473
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1474
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1475
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1476
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1477
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1478
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1479
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1480
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1481
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1482
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1483
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1484
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1485
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1486
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1487
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1488
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1489
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1490
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1491
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1492
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1493
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1494
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1495
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1496
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1497
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1498
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1499
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1500
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1501
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1502
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1503
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1504
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1505
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1506
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1507
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1508
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1509
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1510
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1511
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1512
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1513
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1514
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1515
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1516
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1517
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1518
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1519
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1520
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1521
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1522
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1523
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1524
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1525
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1526
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1527
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1528
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1529
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1530
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1531
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1532
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1533
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1534
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1535
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1536
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1537
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1538
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1539
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1540
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1541
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1542
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1543
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1544
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1545
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1546
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1547
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1548
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1549
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1550
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1551
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1552
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1553
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1554
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1555
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1556
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1557
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1558
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1559
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1560
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1561
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1562
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1563
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1564
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1565
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1566
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1567
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1568
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1569
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1570
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1571
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1572
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1573
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1574
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1575
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1576
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1577
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1578
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1579
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1580
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1581
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1582
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1583
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1584
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1585
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1586
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1587
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1588
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1589
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1590
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1591
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1592
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1593
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1594
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1595
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1596
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1597
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1598
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1599
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1600
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1601
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1602
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1603
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1604
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1605
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1606
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1607
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1608
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1609
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1610
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1611
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1612
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1613
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1614
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1615
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1616
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1617
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1618
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1619
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1620
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1621
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1622
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1623
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1624
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1625
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1626
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1627
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1628
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1629
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1630
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1631
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1632
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1633
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1634
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1635
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1636
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1637
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1638
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1639
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1640
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1641
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1642
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1643
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1644
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1645
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1646
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1647
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1648
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1649
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1650
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1651
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1652
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1653
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1654
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1655
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1656
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1657
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1658
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1659
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1660
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1661
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1662
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1663
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1664
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1665
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1666
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1667
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1668
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1669
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1670
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1671
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1672
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1673
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1674
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1675
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1676
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1677
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1678
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1679
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1680
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1681
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1682
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1683
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1684
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1685
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1686
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1687
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1688
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1689
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1690
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1691
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1692
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1693
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1694
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1695
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1696
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1697
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1698
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1699
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1700
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1701
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1702
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1703
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1704
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1705
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1706
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1707
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1708
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1709
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1710
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1711
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1712
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1713
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1714
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1715
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1716
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1717
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1718
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1719
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1720
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1721
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1722
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1723
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1724
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1725
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1726
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1727
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1728
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1729
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1730
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1731
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1732
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1733
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1734
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1735
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1736
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1737
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1738
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1739
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1740
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1741
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1742
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1743
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1744
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1745
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1746
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1747
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1748
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1749
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1750
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1751
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1752
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1753
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1754
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1755
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1756
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1757
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1758
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1759
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1760
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1761
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1762
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1763
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1764
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1765
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1766
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1767
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1768
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1769
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1770
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1771
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1772
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1773
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1774
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1775
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1776
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1777
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1778
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1779
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1780
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1781
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1782
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1783
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1784
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1785
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1786
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1787
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1788
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1789
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1790
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1791
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1792
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1793
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1794
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1795
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1796
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1797
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1798
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1799
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1800
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1801
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1802
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1803
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1804
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1805
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1806
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1807
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1808
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1809
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1810
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1811
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1812
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1813
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1814
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1815
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1816
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1817
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1818
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1819
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1820
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1821
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1822
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1823
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1824
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1825
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1826
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1827
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1828
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1829
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1830
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1831
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1832
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1833
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1834
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1835
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1836
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1837
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1838
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1839
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1840
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1841
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1842
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1843
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1844
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1845
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1846
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1847
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1848
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1849
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1850
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1851
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1852
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1853
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1854
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1855
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1856
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1857
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1858
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1859
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1860
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1861
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1862
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1863
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1864
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1865
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1866
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1867
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1868
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1869
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1870
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1871
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1872
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1873
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1874
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1875
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1876
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1877
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1878
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1879
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1880
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1881
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1882
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1883
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1884
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1885
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1886
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1887
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1888
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1889
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1890
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1891
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1892
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1893
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1894
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1895
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1896
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1897
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1898
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1899
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1900
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1901
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1902
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1903
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1904
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1905
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1906
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1907
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1908
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1909
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1910
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1911
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1912
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1913
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1914
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1915
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1916
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1917
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1918
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1919
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1920
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1921
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1922
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1923
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1924
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1925
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1926
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1927
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1928
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1929
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1930
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1931
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1932
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1933
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1934
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1935
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1936
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1937
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1938
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1939
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1940
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1941
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1942
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1943
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1944
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1945
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1946
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1947
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1948
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1949
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1950
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1951
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1952
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1953
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1954
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1955
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1956
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1957
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1958
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1959
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1960
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1961
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1962
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1963
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1964
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1965
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1966
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1967
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1968
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1969
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1970
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1971
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1972
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1973
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1974
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1975
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1976
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1977
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1978
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1979
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1980
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1981
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1982
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1983
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1984
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1985
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1986
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1987
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1988
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1989
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1990
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1991
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1992
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1993
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1994
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1995
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1996
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1997
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1998
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 1999
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 2000
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 2001
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 2002
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        -- instruction 2003
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);
        
        uart_buffer_write <= '1';
        uart_data_in <= x"00";
        
        wait until rising_edge(clk_sig);
        uart_buffer_write <= '0';
        
        wait until uart_tx_buf_pres = '0';
        wait until rising_edge(clk_sig);

        
        wait for 50000ms;
    end process simulate;
end Behavioral;
